module CPU_module (

);
// Do not use me (yet)

endmodule
